library verilog;
use verilog.vl_types.all;
entity UART_5_vlg_vec_tst is
end UART_5_vlg_vec_tst;
